`define CPU_CYCLE     10.0 // 100Mhz
`define MAX           10000000//207569
