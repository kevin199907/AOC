module control(
		input clk,
		input rst,
		output logic[13:0]A,
		output logic WM_OE,
		input  logic[31:0]DO,
		input  logic fifo_WREADY_row    [15:0][15:0],
		output logic fifo_WVALID_row    [15:0][15:0],
		output logic [7:0]    in_row    [15:0][15:0],
		output logic [6:0]    state
);

integer i;
integer j;
always@(posedge clk)begin:sadasd
	if(rst)begin
	A<=0;
	 WM_OE<=0;

	state<=0;
			end
		

	else if(state<68)begin
	WM_OE<=1;
	A<=A+1;
	state<=state+1;
	end
	//else if(state==68)begin
	//state<=0;
	//WM_OE<=1;
	//end
	
	else begin
	WM_OE<=0;
	A<=A;
	for(i=0;i<16;i=i+1)begin
		for(j=0;j<16;j=j+1)
			fifo_WVALID_row[i][j]<=1'd0;
			end
	state<=state;
	end

end

always@(posedge clk)begin
	case(state)
//=============pointwise1============================================================

	7'd1:begin	
	 in_row[0][0]<=DO[7:0];
	 in_row[0][1]<=DO[15:8];
	 in_row[0][2]<=DO[23:16];
	 in_row[0][3]<=DO[31:24];
	fifo_WVALID_row[0][0]<=1'd1;
    fifo_WVALID_row[0][1]<=1'd1;
    fifo_WVALID_row[0][2]<=1'd1;
    fifo_WVALID_row[0][3]<=1'd1;			
	end
	7'd2:begin

	fifo_WVALID_row[0][0]<=1'd0;
    fifo_WVALID_row[0][1]<=1'd0;
    fifo_WVALID_row[0][2]<=1'd0;
    fifo_WVALID_row[0][3]<=1'd0;
	
	fifo_WVALID_row[0][7]<=1'd1;
	fifo_WVALID_row[0][6]<=1'd1;
	fifo_WVALID_row[0][5]<=1'd1;
	fifo_WVALID_row[0][4]<=1'd1;
	in_row[0][4]<=DO[7:0];
	in_row[0][5]<=DO[15:8];
	in_row[0][6]<=DO[23:16];
	in_row[0][7]<=DO[31:24];
	end	
	7'd3:begin
	
	fifo_WVALID_row[0][4]<=1'd0;
	fifo_WVALID_row[0][5]<=1'd0;
	fifo_WVALID_row[0][6]<=1'd0;
	fifo_WVALID_row[0][7]<=1'd0;
	
			 in_row[1][0]<=DO[7:0];
			 in_row[1][1]<=DO[15:8];
			 in_row[1][2]<=DO[23:16];
			 in_row[1][3]<=DO[31:24];
	fifo_WVALID_row[1][0]<=1'd1;
    fifo_WVALID_row[1][1]<=1'd1;
    fifo_WVALID_row[1][2]<=1'd1;
    fifo_WVALID_row[1][3]<=1'd1;	
	end	
	7'd4:begin//////////////////////////////////////////////////////
	fifo_WVALID_row[1][0]<=1'd0;
    fifo_WVALID_row[1][1]<=1'd0;
    fifo_WVALID_row[1][2]<=1'd0;
    fifo_WVALID_row[1][3]<=1'd0;
	
			 in_row[1][4]<=DO[7:0];
			 in_row[1][5]<=DO[15:8];
			 in_row[1][6]<=DO[23:16];
			 in_row[1][7]<=DO[31:24];
	fifo_WVALID_row[1][4]<=1'd1;
    fifo_WVALID_row[1][5]<=1'd1;
    fifo_WVALID_row[1][6]<=1'd1;
    fifo_WVALID_row[1][7]<=1'd1;		
	end	
	7'd5:begin
	fifo_WVALID_row[1][4]<=1'd0;
    fifo_WVALID_row[1][5]<=1'd0;
    fifo_WVALID_row[1][6]<=1'd0;
    fifo_WVALID_row[1][7]<=1'd0;
	
			 in_row[2][0]<=DO[7:0];
			 in_row[2][1]<=DO[15:8];
			 in_row[2][2]<=DO[23:16];
			 in_row[2][3]<=DO[31:24];
	fifo_WVALID_row[2][0]<=1'd1;
    fifo_WVALID_row[2][1]<=1'd1;
    fifo_WVALID_row[2][2]<=1'd1;
    fifo_WVALID_row[2][3]<=1'd1;		
	end	
	7'd6:begin
	fifo_WVALID_row[2][0]<=1'd0;
    fifo_WVALID_row[2][1]<=1'd0;
    fifo_WVALID_row[2][2]<=1'd0;
    fifo_WVALID_row[2][3]<=1'd0;
			 in_row[2][4]<=DO[7:0];
			 in_row[2][5]<=DO[15:8];
			 in_row[2][6]<=DO[23:16];
			 in_row[2][7]<=DO[31:24];
	fifo_WVALID_row[2][4]<=1'd1;
    fifo_WVALID_row[2][5]<=1'd1;
    fifo_WVALID_row[2][6]<=1'd1;
    fifo_WVALID_row[2][7]<=1'd1;	
	end	
	7'd7:begin
	fifo_WVALID_row[2][4]<=1'd0;
    fifo_WVALID_row[2][5]<=1'd0;
    fifo_WVALID_row[2][6]<=1'd0;
    fifo_WVALID_row[2][7]<=1'd0;
	in_row[3][0]<=DO[7:0];
	in_row[3][1]<=DO[15:8];
	in_row[3][2]<=DO[23:16];
	in_row[3][3]<=DO[31:24];
	fifo_WVALID_row[3][0]<=1'd1;
    fifo_WVALID_row[3][1]<=1'd1;
    fifo_WVALID_row[3][2]<=1'd1;
    fifo_WVALID_row[3][3]<=1'd1;	
	end	
	7'd8:begin
	fifo_WVALID_row[3][0]<=1'd0;
    fifo_WVALID_row[3][1]<=1'd0;
    fifo_WVALID_row[3][2]<=1'd0;
    fifo_WVALID_row[3][3]<=1'd0;	
	in_row[3][4]<=DO[7:0];
	in_row[3][5]<=DO[15:8];
	in_row[3][6]<=DO[23:16];
	in_row[3][7]<=DO[31:24];
	fifo_WVALID_row[3][4]<=1'd1;
    fifo_WVALID_row[3][5]<=1'd1;
    fifo_WVALID_row[3][6]<=1'd1;
    fifo_WVALID_row[3][7]<=1'd1;		
	end	
	7'd9:begin
	fifo_WVALID_row[3][4]<=1'd0;
    fifo_WVALID_row[3][5]<=1'd0;
    fifo_WVALID_row[3][6]<=1'd0;
    fifo_WVALID_row[3][7]<=1'd0;
	in_row[4][0]<=DO[7:0];
	in_row[4][1]<=DO[15:8];
	in_row[4][2]<=DO[23:16];
	in_row[4][3]<=DO[31:24];
	fifo_WVALID_row[4][0]<=1'd1;
    fifo_WVALID_row[4][1]<=1'd1;
    fifo_WVALID_row[4][2]<=1'd1;
    fifo_WVALID_row[4][3]<=1'd1;	
	end	
	7'd10:begin//////////////////
	fifo_WVALID_row[4][0]<=1'd0;
    fifo_WVALID_row[4][1]<=1'd0;
    fifo_WVALID_row[4][2]<=1'd0;
    fifo_WVALID_row[4][3]<=1'd0;
	in_row[4][4]<=DO[7:0];
	in_row[4][5]<=DO[15:8];
	in_row[4][6]<=DO[23:16];
	in_row[4][7]<=DO[31:24];
	fifo_WVALID_row[4][4]<=1'd1;
    fifo_WVALID_row[4][5]<=1'd1;
    fifo_WVALID_row[4][6]<=1'd1;
    fifo_WVALID_row[4][7]<=1'd1;	
	end	
	7'd11:begin
	fifo_WVALID_row[4][4]<=1'd0;
    fifo_WVALID_row[4][5]<=1'd0;
    fifo_WVALID_row[4][6]<=1'd0;
    fifo_WVALID_row[4][7]<=1'd0;	
	in_row[5][0]<=DO[7:0];
	in_row[5][1]<=DO[15:8];
	in_row[5][2]<=DO[23:16];
	in_row[5][3]<=DO[31:24];
	fifo_WVALID_row[5][0]<=1'd1;
    fifo_WVALID_row[5][1]<=1'd1;
    fifo_WVALID_row[5][2]<=1'd1;
    fifo_WVALID_row[5][3]<=1'd1;		
	end	
	7'd12:begin
	fifo_WVALID_row[5][0]<=1'd0;
    fifo_WVALID_row[5][1]<=1'd0;
    fifo_WVALID_row[5][2]<=1'd0;
    fifo_WVALID_row[5][3]<=1'd0;
	in_row[5][4]<=DO[7:0];
	in_row[5][5]<=DO[15:8];
	in_row[5][6]<=DO[23:16];
	in_row[5][7]<=DO[31:24];
	fifo_WVALID_row[5][4]<=1'd1;
    fifo_WVALID_row[5][5]<=1'd1;
    fifo_WVALID_row[5][6]<=1'd1;
    fifo_WVALID_row[5][7]<=1'd1;	
	end	
	7'd13:begin
	fifo_WVALID_row[5][4]<=1'd0;
    fifo_WVALID_row[5][5]<=1'd0;
    fifo_WVALID_row[5][6]<=1'd0;
    fifo_WVALID_row[5][7]<=1'd0;
	in_row[6][0]<=DO[7:0];
	in_row[6][1]<=DO[15:8];
	in_row[6][2]<=DO[23:16];
	in_row[6][3]<=DO[31:24];
	fifo_WVALID_row[6][0]<=1'd1;
    fifo_WVALID_row[6][1]<=1'd1;
    fifo_WVALID_row[6][2]<=1'd1;
    fifo_WVALID_row[6][3]<=1'd1;	
	end	
	7'd14:begin
	fifo_WVALID_row[6][0]<=1'd0;
    fifo_WVALID_row[6][1]<=1'd0;
    fifo_WVALID_row[6][2]<=1'd0;
    fifo_WVALID_row[6][3]<=1'd0;	
	in_row[6][4]<=DO[7:0];
	in_row[6][5]<=DO[15:8];
	in_row[6][6]<=DO[23:16];
	in_row[6][7]<=DO[31:24];
	fifo_WVALID_row[6][4]<=1'd1;
    fifo_WVALID_row[6][5]<=1'd1;
    fifo_WVALID_row[6][6]<=1'd1;
    fifo_WVALID_row[6][7]<=1'd1;		
	end		
	7'd15:begin
	fifo_WVALID_row[6][4]<=1'd0;
    fifo_WVALID_row[6][5]<=1'd0;
    fifo_WVALID_row[6][6]<=1'd0;
    fifo_WVALID_row[6][7]<=1'd0;
	in_row[7][0]<=DO[7:0];
	in_row[7][1]<=DO[15:8];
	in_row[7][2]<=DO[23:16];
	in_row[7][3]<=DO[31:24];
	fifo_WVALID_row[7][0]<=1'd1;
    fifo_WVALID_row[7][1]<=1'd1;
    fifo_WVALID_row[7][2]<=1'd1;
    fifo_WVALID_row[7][3]<=1'd1;	
	end	
	7'd16:begin
	fifo_WVALID_row[7][0]<=1'd0;
    fifo_WVALID_row[7][1]<=1'd0;
    fifo_WVALID_row[7][2]<=1'd0;
    fifo_WVALID_row[7][3]<=1'd0;	
	in_row[7][4]<=DO[7:0];
	in_row[7][5]<=DO[15:8];
	in_row[7][6]<=DO[23:16];
	in_row[7][7]<=DO[31:24];
	fifo_WVALID_row[7][4]<=1'd1;
    fifo_WVALID_row[7][5]<=1'd1;
    fifo_WVALID_row[7][6]<=1'd1;
    fifo_WVALID_row[7][7]<=1'd1;	
	end	
//=============pointwise1============================================================	
//=============depthwise1============================================================	
	7'd17:begin
	fifo_WVALID_row[7][4]<=1'd0;
    fifo_WVALID_row[7][5]<=1'd0;
    fifo_WVALID_row[7][6]<=1'd0;
    fifo_WVALID_row[7][7]<=1'd0;
	in_row[2][0]<=DO[7:0];
	in_row[2][1]<=DO[15:8];
	in_row[2][2]<=DO[23:16];
	in_row[1][0]<=DO[31:24];
	fifo_WVALID_row[2][0]<=1'd1;
    fifo_WVALID_row[2][1]<=1'd1;
    fifo_WVALID_row[2][2]<=1'd1;
    fifo_WVALID_row[1][0]<=1'd1;	
	end	
	7'd18:begin
	fifo_WVALID_row[2][0]<=1'd0;
    fifo_WVALID_row[2][1]<=1'd0;
    fifo_WVALID_row[2][2]<=1'd0;
    fifo_WVALID_row[1][0]<=1'd0;
	in_row[1][1]<=DO[7:0];
	in_row[1][2]<=DO[15:8];
	in_row[0][0]<=DO[23:16];
	in_row[0][1]<=DO[31:24];
	fifo_WVALID_row[1][1]<=1'd1;
    fifo_WVALID_row[1][2]<=1'd1;
    fifo_WVALID_row[0][0]<=1'd1;
    fifo_WVALID_row[0][1]<=1'd1;	
	end	
	7'd19:begin
	fifo_WVALID_row[1][1]<=1'd0;
    fifo_WVALID_row[1][2]<=1'd0;
    fifo_WVALID_row[0][0]<=1'd0;
    fifo_WVALID_row[0][1]<=1'd0;		
	in_row[0][2]<=DO[7:0];
	in_row[5][3]<=DO[15:8];
	in_row[5][4]<=DO[23:16];
	in_row[5][5]<=DO[31:24];
	fifo_WVALID_row[0][2]<=1'd1;
    fifo_WVALID_row[5][3]<=1'd1;
    fifo_WVALID_row[5][4]<=1'd1;
    fifo_WVALID_row[5][5]<=1'd1;		
	end	
	7'd20:begin
	fifo_WVALID_row[0][2]<=1'd0;
    fifo_WVALID_row[5][3]<=1'd0;
    fifo_WVALID_row[5][4]<=1'd0;
    fifo_WVALID_row[5][5]<=1'd0;
	in_row[4][3]<=DO[7:0];
	in_row[4][4]<=DO[15:8];
	in_row[4][5]<=DO[23:16];
	in_row[3][3]<=DO[31:24];
	fifo_WVALID_row[4][3]<=1'd1;
    fifo_WVALID_row[4][4]<=1'd1;
    fifo_WVALID_row[4][5]<=1'd1;
    fifo_WVALID_row[3][3]<=1'd1;	
	end	
	7'd21:begin
	fifo_WVALID_row[4][3]<=1'd0;
    fifo_WVALID_row[4][4]<=1'd0;
    fifo_WVALID_row[4][5]<=1'd0;
    fifo_WVALID_row[3][3]<=1'd0;
	in_row[3][4]<=DO[7:0];
	in_row[3][5]<=DO[15:8];	      
	in_row[8][6]<=DO[23:16];
	in_row[8][7]<=DO[31:24];
	fifo_WVALID_row[3][4]<=1'd1;
    fifo_WVALID_row[3][5]<=1'd1;
    fifo_WVALID_row[8][6]<=1'd1;
    fifo_WVALID_row[8][7]<=1'd1;	
	end	
	7'd22:begin
	fifo_WVALID_row[3][4]<=1'd0;
    fifo_WVALID_row[3][5]<=1'd0;
    fifo_WVALID_row[8][6]<=1'd0;
    fifo_WVALID_row[8][7]<=1'd0;
	in_row[8][8]<=DO[7:0];
	in_row[7][6]<=DO[15:8];
	in_row[7][7]<=DO[23:16];
	in_row[7][8]<=DO[31:24];
	fifo_WVALID_row[8][8]<=1'd1;
    fifo_WVALID_row[7][6]<=1'd1;
    fifo_WVALID_row[7][7]<=1'd1;
    fifo_WVALID_row[7][8]<=1'd1;	
	end	
	7'd23:begin
	fifo_WVALID_row[8][8]<=1'd0;
    fifo_WVALID_row[7][6]<=1'd0;
    fifo_WVALID_row[7][7]<=1'd0;
    fifo_WVALID_row[7][8]<=1'd0;
	in_row[6][6] <=DO[7:0];
	in_row[6][7] <=DO[15:8];
	in_row[6][8] <=DO[23:16];
	in_row[11][9]<=DO[31:24];
	fifo_WVALID_row[6][6] <=1'd1;
    fifo_WVALID_row[6][7] <=1'd1;
    fifo_WVALID_row[6][8] <=1'd1;
    fifo_WVALID_row[11][9]<=1'd1;	
	
	end	
	7'd24:begin
	fifo_WVALID_row[6][6] <=1'd0;
    fifo_WVALID_row[6][7] <=1'd0;
    fifo_WVALID_row[6][8] <= 1'd0;
    fifo_WVALID_row[11][9]<=1'd0;	
	in_row[11][10]<=DO[7:0];
	in_row[11][11]<=DO[15:8];
	in_row[10][9] <=DO[23:16];
	in_row[10][10]<=DO[31:24];
	fifo_WVALID_row[11][10]<=1'd1;
    fifo_WVALID_row[11][11]<=1'd1;
    fifo_WVALID_row[10][9] <= 1'd1;
    fifo_WVALID_row[10][10]<=1'd1;	
	end	
	7'd25:begin
	fifo_WVALID_row[11][10]<=1'd0;
    fifo_WVALID_row[11][11]<=1'd0;
    fifo_WVALID_row[10][9] <=1'd0;
    fifo_WVALID_row[10][10]<=1'd0;	
	in_row[10][11]<=DO[7:0];
	in_row[9][9]  <=DO[15:8];
	in_row[9][10] <=DO[23:16];
	in_row[9][11] <=DO[31:24];	
	fifo_WVALID_row[10][11]<=1'd1;
    fifo_WVALID_row[9][9]  <=1'd1;
    fifo_WVALID_row[9][10] <= 1'd1;
    fifo_WVALID_row[9][11] <=1'd1;	
	end	
	7'd26:begin
	fifo_WVALID_row[10][11]<=1'd0;
    fifo_WVALID_row[9][9]  <=1'd0;
    fifo_WVALID_row[9][10] <=1'd0;
    fifo_WVALID_row[9][11] <=1'd0;	
	in_row[14][12]<=DO[7:0];
	in_row[14][13]<=DO[15:8];
	in_row[14][14]<=DO[23:16];
	in_row[13][12]<=DO[31:24];	
	fifo_WVALID_row[14][12]<=1'd1;
    fifo_WVALID_row[14][13]<=1'd1;
    fifo_WVALID_row[14][14]<= 1'd1;
    fifo_WVALID_row[13][12]<=1'd1;	
	end	
	7'd27:begin
	fifo_WVALID_row[14][12]<=1'd0;
    fifo_WVALID_row[14][13]<=1'd0;
    fifo_WVALID_row[14][14]<=1'd0;
    fifo_WVALID_row[13][12]<=1'd0;	
	in_row[13][13]<=DO[7:0];
	in_row[13][14]<=DO[15:8];
	in_row[12][12]<=DO[23:16];
	in_row[12][13]<=DO[31:24];
	fifo_WVALID_row[13][13]<=1'd1;
    fifo_WVALID_row[13][14]<=1'd1;
    fifo_WVALID_row[12][12]<=1'd1;
    fifo_WVALID_row[12][13]<=1'd1;		
	end	
	7'd28:begin
	fifo_WVALID_row[13][13]<=1'd0;
    fifo_WVALID_row[13][14]<=1'd0;
    fifo_WVALID_row[12][12]<=1'd0;
    fifo_WVALID_row[12][13]<=1'd0;
	in_row[12][14]<=DO[7:0];
//=============depthwise1============================================================
//=============depthwise2============================================================
	in_row[2][0]<=DO[15:8];
	in_row[2][1]<=DO[23:16];
	in_row[2][2]<=DO[31:24];
	fifo_WVALID_row[12][14]<=1'd1;
    fifo_WVALID_row[2][0]<=1'd1;
    fifo_WVALID_row[2][1]<=1'd1;
    fifo_WVALID_row[2][2]<=1'd1;
	end	
	7'd29:begin
	fifo_WVALID_row[12][14]<=1'd0;
    fifo_WVALID_row[2][0]<=1'd0;
    fifo_WVALID_row[2][1]<=1'd0;
    fifo_WVALID_row[2][2]<=1'd0;
	in_row[1][0]<=DO[7:0];
	in_row[1][1]<=DO[15:8];
	in_row[1][2]<=DO[23:16];
	in_row[0][0]<=DO[31:24];
	fifo_WVALID_row[1][0]<=1'd1;
    fifo_WVALID_row[1][1]<=1'd1;
    fifo_WVALID_row[1][2]<=1'd1;
    fifo_WVALID_row[0][0]<=1'd1;	
	end	
	7'd30:begin
	fifo_WVALID_row[1][0]<=1'd0;
    fifo_WVALID_row[1][1]<=1'd0;
    fifo_WVALID_row[1][2]<=1'd0;
    fifo_WVALID_row[0][0]<=1'd0;	
	in_row[0][1]<=DO[7:0];
	in_row[0][2]<=DO[15:8];
	in_row[5][3]<=DO[23:16];
	in_row[5][4]<=DO[31:24];
	fifo_WVALID_row[0][1]<=1'd1;
    fifo_WVALID_row[0][2]<=1'd1;
    fifo_WVALID_row[5][3]<=1'd1;
    fifo_WVALID_row[5][4]<=1'd1;		
	end
	7'd31:begin////////////////////
	fifo_WVALID_row[0][1]<=1'd0;
    fifo_WVALID_row[0][2]<=1'd0;
    fifo_WVALID_row[5][3]<=1'd0;
    fifo_WVALID_row[5][4]<=1'd0;
	in_row[5][5]<=DO[7:0];
	in_row[4][3]<=DO[15:8];
	in_row[4][4]<=DO[23:16];
	in_row[4][5]<=DO[31:24];
	fifo_WVALID_row[5][5]<=1'd1;
    fifo_WVALID_row[4][3]<=1'd1;
    fifo_WVALID_row[4][4]<=1'd1;
    fifo_WVALID_row[4][5]<=1'd1;	
	end		
	7'd32:begin
	fifo_WVALID_row[5][5]<=1'd0;
    fifo_WVALID_row[4][3]<=1'd0;
    fifo_WVALID_row[4][4]<=1'd0;
    fifo_WVALID_row[4][5]<=1'd0;
	in_row[3][3]<=DO[7:0];
	in_row[3][4]<=DO[15:8];
	in_row[3][5]<=DO[23:16];
	in_row[8][6]<=DO[31:24];
	fifo_WVALID_row[3][3]<=1'd1;
    fifo_WVALID_row[3][4]<=1'd1;
    fifo_WVALID_row[3][5]<=1'd1;
    fifo_WVALID_row[8][6]<=1'd1;	
	end	
	7'd33:begin
	fifo_WVALID_row[3][3]<=1'd0;
    fifo_WVALID_row[3][4]<=1'd0;
    fifo_WVALID_row[3][5]<=1'd0;
    fifo_WVALID_row[8][6]<=1'd0;	
	in_row[8][7]<=DO[7:0];
	in_row[8][8]<=DO[15:8];
	in_row[7][6]<=DO[23:16];
	in_row[7][7]<=DO[31:24];
	fifo_WVALID_row[8][7]<=1'd1;
    fifo_WVALID_row[8][8]<=1'd1;
    fifo_WVALID_row[7][6]<=1'd1;
    fifo_WVALID_row[7][7]<=1'd1;		
	end	
	7'd34:begin
	fifo_WVALID_row[8][7]<=1'd0;
    fifo_WVALID_row[8][8]<=1'd0;
    fifo_WVALID_row[7][6]<=1'd0;
    fifo_WVALID_row[7][7]<=1'd0;
	in_row[7][8]<=DO[7:0];
	in_row[6][6]<=DO[15:8];
	in_row[6][7]<=DO[23:16];
	in_row[6][8]<=DO[31:24];
	fifo_WVALID_row[7][8]<=1'd1;
    fifo_WVALID_row[6][6]<=1'd1;
    fifo_WVALID_row[6][7]<=1'd1;
    fifo_WVALID_row[6][8]<=1'd1;	
	end		
//=============depthwise2============================================================				
//=============pointwise2============================================================	
	7'd35:begin
	fifo_WVALID_row[7][8]<=1'd0;
    fifo_WVALID_row[6][6]<=1'd0;
    fifo_WVALID_row[6][7]<=1'd0;
    fifo_WVALID_row[6][8]<=1'd0;	
	in_row[0][0]<=DO[7:0];
	in_row[0][1]<=DO[15:8];
	in_row[0][2]<=DO[23:16];
	in_row[0][3]<=DO[31:24];
	fifo_WVALID_row[0][0]<=1'd1;
    fifo_WVALID_row[0][1]<=1'd1;
    fifo_WVALID_row[0][2]<=1'd1;
    fifo_WVALID_row[0][3]<=1'd1;		
	end
	7'd36:begin
	fifo_WVALID_row[0][0]<=1'd0;
	fifo_WVALID_row[0][1]<=1'd0;
	fifo_WVALID_row[0][2]<=1'd0;
	fifo_WVALID_row[0][3]<=1'd0;
	in_row[0][4]<=DO[7:0];
	in_row[0][5]<=DO[15:8];
	in_row[0][6]<=DO[23:16];
	in_row[0][7]<=DO[31:24];
	fifo_WVALID_row[0][4]<=1'd1;
    fifo_WVALID_row[0][5]<=1'd1;
    fifo_WVALID_row[0][6]<=1'd1;
    fifo_WVALID_row[0][7]<=1'd1;
	end	
	7'd37:begin
	fifo_WVALID_row[0][4]<=1'd0;
    fifo_WVALID_row[0][5]<=1'd0;
    fifo_WVALID_row[0][6]<=1'd0;
    fifo_WVALID_row[0][7]<=1'd0;	
	in_row[1][0]<=DO[7:0];
	in_row[1][1]<=DO[15:8];
	in_row[1][2]<=DO[23:16];
	in_row[1][3]<=DO[31:24];
	fifo_WVALID_row[1][0]<=1'd1;
    fifo_WVALID_row[1][1]<=1'd1;
    fifo_WVALID_row[1][2]<=1'd1;
    fifo_WVALID_row[1][3]<=1'd1;
	end	
	7'd38:begin
	fifo_WVALID_row[1][0]<=1'd0;
    fifo_WVALID_row[1][1]<=1'd0;
    fifo_WVALID_row[1][2]<=1'd0;
    fifo_WVALID_row[1][3]<=1'd0;	
	in_row[1][4]<=DO[7:0];
	in_row[1][5]<=DO[15:8];
	in_row[1][6]<=DO[23:16];
	in_row[1][7]<=DO[31:24];
	fifo_WVALID_row[1][4]<=1'd1;
    fifo_WVALID_row[1][5]<=1'd1;
    fifo_WVALID_row[1][6]<=1'd1;
    fifo_WVALID_row[1][7]<=1'd1;
	end	
	7'd39:begin
	fifo_WVALID_row[1][4]<=1'd0;
    fifo_WVALID_row[1][5]<=1'd0;
    fifo_WVALID_row[1][6]<=1'd0;
    fifo_WVALID_row[1][7]<=1'd0;	
	in_row[2][0]<=DO[7:0];
	in_row[2][1]<=DO[15:8];
	in_row[2][2]<=DO[23:16];
	in_row[2][3]<=DO[31:24];
	fifo_WVALID_row[2][0]<=1'd1;
    fifo_WVALID_row[2][1]<=1'd1;
    fifo_WVALID_row[2][2]<=1'd1;
    fifo_WVALID_row[2][3]<=1'd1;	
	end	
	7'd40:begin
	fifo_WVALID_row[2][0]<=1'd0;
    fifo_WVALID_row[2][1]<=1'd0;
    fifo_WVALID_row[2][2]<=1'd0;
    fifo_WVALID_row[2][3]<=1'd0;
	in_row[2][4]<=DO[7:0];
	in_row[2][5]<=DO[15:8];
	in_row[2][6]<=DO[23:16];
	in_row[2][7]<=DO[31:24];
	fifo_WVALID_row[2][4]<=1'd1;
    fifo_WVALID_row[2][5]<=1'd1;
    fifo_WVALID_row[2][6]<=1'd1;
    fifo_WVALID_row[2][7]<=1'd1;	
	end	
	7'd41:begin
	fifo_WVALID_row[2][4]<=1'd0;
    fifo_WVALID_row[2][5]<=1'd0;
    fifo_WVALID_row[2][6]<=1'd0;
    fifo_WVALID_row[2][7]<=1'd0;
	in_row[3][0]<=DO[7:0];
	in_row[3][1]<=DO[15:8];
	in_row[3][2]<=DO[23:16];
	in_row[3][3]<=DO[31:24];
	fifo_WVALID_row[3][0]<=1'd1;
    fifo_WVALID_row[3][1]<=1'd1;
    fifo_WVALID_row[3][2]<=1'd1;
    fifo_WVALID_row[3][3]<=1'd1;	
	end	
	7'd42:begin
	fifo_WVALID_row[3][0]<=1'd0;
    fifo_WVALID_row[3][1]<=1'd0;
    fifo_WVALID_row[3][2]<=1'd0;
    fifo_WVALID_row[3][3]<=1'd0;	
	in_row[3][4]<=DO[7:0];
	in_row[3][5]<=DO[15:8];
	in_row[3][6]<=DO[23:16];
	in_row[3][7]<=DO[31:24];
	fifo_WVALID_row[3][4]<=1'd1;
    fifo_WVALID_row[3][5]<=1'd1;
    fifo_WVALID_row[3][6]<=1'd1;
    fifo_WVALID_row[3][7]<=1'd1;		
	end	
	7'd43:begin
	fifo_WVALID_row[3][4]<=1'd0;
    fifo_WVALID_row[3][5]<=1'd0;
    fifo_WVALID_row[3][6]<=1'd0;
    fifo_WVALID_row[3][7]<=1'd0;
	in_row[4][0]<=DO[7:0];
	in_row[4][1]<=DO[15:8];
	in_row[4][2]<=DO[23:16];
	in_row[4][3]<=DO[31:24];
	fifo_WVALID_row[4][0]<=1'd1;
    fifo_WVALID_row[4][1]<=1'd1;
    fifo_WVALID_row[4][2]<=1'd1;
    fifo_WVALID_row[4][3]<=1'd1;	
	end	
	7'd44:begin
	fifo_WVALID_row[4][0]<=1'd0;
    fifo_WVALID_row[4][1]<=1'd0;
    fifo_WVALID_row[4][2]<=1'd0;
    fifo_WVALID_row[4][3]<=1'd0;
	in_row[4][4]<=DO[7:0];
	in_row[4][5]<=DO[15:8];
	in_row[4][6]<=DO[23:16];
	in_row[4][7]<=DO[31:24];
	fifo_WVALID_row[4][4]<=1'd1;
    fifo_WVALID_row[4][5]<=1'd1;
    fifo_WVALID_row[4][6]<=1'd1;
    fifo_WVALID_row[4][7]<=1'd1;	
	end	
	7'd45:begin
	fifo_WVALID_row[4][4]<=1'd0;
    fifo_WVALID_row[4][5]<=1'd0;
    fifo_WVALID_row[4][6]<=1'd0;
    fifo_WVALID_row[4][7]<=1'd0;	
	in_row[5][0]<=DO[7:0];
	in_row[5][1]<=DO[15:8];
	in_row[5][2]<=DO[23:16];
	in_row[5][3]<=DO[31:24];
	fifo_WVALID_row[5][0]<=1'd1;
    fifo_WVALID_row[5][1]<=1'd1;
    fifo_WVALID_row[5][2]<=1'd1;
    fifo_WVALID_row[5][3]<=1'd1;	
	end	
	7'd46:begin
	fifo_WVALID_row[5][0]<=1'd0;
    fifo_WVALID_row[5][1]<=1'd0;
    fifo_WVALID_row[5][2]<=1'd0;
    fifo_WVALID_row[5][3]<=1'd0;
	in_row[5][4]<=DO[7:0];
	in_row[5][5]<=DO[15:8];
	in_row[5][6]<=DO[23:16];
	in_row[5][7]<=DO[31:24];
	fifo_WVALID_row[5][4]<=1'd1;
    fifo_WVALID_row[5][5]<=1'd1;
    fifo_WVALID_row[5][6]<=1'd1;
    fifo_WVALID_row[5][7]<=1'd1;
	end	
	7'd47:begin
	fifo_WVALID_row[5][4]<=1'd0;
    fifo_WVALID_row[5][5]<=1'd0;
    fifo_WVALID_row[5][6]<=1'd0;
    fifo_WVALID_row[5][7]<=1'd0;
	in_row[6][0]<=DO[7:0];
	in_row[6][1]<=DO[15:8];
	in_row[6][2]<=DO[23:16];
	in_row[6][3]<=DO[31:24];
	fifo_WVALID_row[6][0]<=1'd1;
    fifo_WVALID_row[6][1]<=1'd1;
    fifo_WVALID_row[6][2]<=1'd1;
    fifo_WVALID_row[6][3]<=1'd1;	
	end	
	7'd48:begin///////////////////////////////////////////////////////
	fifo_WVALID_row[6][0]<=1'd0;
    fifo_WVALID_row[6][1]<=1'd0;
    fifo_WVALID_row[6][2]<=1'd0;
    fifo_WVALID_row[6][3]<=1'd0;	
	in_row[6][4]<=DO[7:0];
	in_row[6][5]<=DO[15:8];
	in_row[6][6]<=DO[23:16];
	in_row[6][7]<=DO[31:24];
	fifo_WVALID_row[6][4]<=1'd1;
    fifo_WVALID_row[6][5]<=1'd1;
    fifo_WVALID_row[6][6]<=1'd1;
    fifo_WVALID_row[6][7]<=1'd1;
	end		
	7'd49:begin
	fifo_WVALID_row[6][4]<=1'd0;
    fifo_WVALID_row[6][5]<=1'd0;
    fifo_WVALID_row[6][6]<=1'd0;
    fifo_WVALID_row[6][7]<=1'd0;
	in_row[7][0]<=DO[7:0];
	in_row[7][1]<=DO[15:8];
	in_row[7][2]<=DO[23:16];
	in_row[7][3]<=DO[31:24];
	fifo_WVALID_row[7][0]<=1'd1;
    fifo_WVALID_row[7][1]<=1'd1;
    fifo_WVALID_row[7][2]<=1'd1;
    fifo_WVALID_row[7][3]<=1'd1;
	end	
	7'd50:begin
	fifo_WVALID_row[7][0]<=1'd0;
    fifo_WVALID_row[7][1]<=1'd0;
    fifo_WVALID_row[7][2]<=1'd0;
    fifo_WVALID_row[7][3]<=1'd0;	
			 in_row[7][4]<=DO[7:0];
			 in_row[7][5]<=DO[15:8];
			 in_row[7][6]<=DO[23:16];
			 in_row[7][7]<=DO[31:24];
	fifo_WVALID_row[7][4]<=1'd1;
    fifo_WVALID_row[7][5]<=1'd1;
    fifo_WVALID_row[7][6]<=1'd1;
    fifo_WVALID_row[7][7]<=1'd1;		
	end	
	7'd51:begin
	fifo_WVALID_row[7][4]<=1'd0;
    fifo_WVALID_row[7][5]<=1'd0;
    fifo_WVALID_row[7][6]<=1'd0;
    fifo_WVALID_row[7][7]<=1'd0;	
	in_row[8][0]<=DO[7:0];
	in_row[8][1]<=DO[15:8];
	in_row[8][2]<=DO[23:16];
	in_row[8][3]<=DO[31:24];
	fifo_WVALID_row[8][0]<=1'd1;
    fifo_WVALID_row[8][1]<=1'd1;
    fifo_WVALID_row[8][2]<=1'd1;
    fifo_WVALID_row[8][3]<=1'd1;		
	end
	7'd52:begin
	fifo_WVALID_row[8][0]<=1'd0;
    fifo_WVALID_row[8][1]<=1'd0;
    fifo_WVALID_row[8][2]<=1'd0;
    fifo_WVALID_row[8][3]<=1'd0;	
	in_row[8][4]<=DO[7:0];
	in_row[8][5]<=DO[15:8];
	in_row[8][6]<=DO[23:16];
	in_row[8][7]<=DO[31:24];
	fifo_WVALID_row[8][4]<=1'd1;
    fifo_WVALID_row[8][5]<=1'd1;
    fifo_WVALID_row[8][6]<=1'd1;
    fifo_WVALID_row[8][7]<=1'd1;		
	end	
	7'd53:begin
	fifo_WVALID_row[8][4]<=1'd0;
    fifo_WVALID_row[8][5]<=1'd0;
    fifo_WVALID_row[8][6]<=1'd0;
    fifo_WVALID_row[8][7]<=1'd0;
	in_row[9][0]<=DO[7:0];
	in_row[9][1]<=DO[15:8];
	in_row[9][2]<=DO[23:16];
	in_row[9][3]<=DO[31:24];
	fifo_WVALID_row[9][0]<=1'd1;
    fifo_WVALID_row[9][1]<=1'd1;
    fifo_WVALID_row[9][2]<=1'd1;
    fifo_WVALID_row[9][3]<=1'd1;	
	end	
	7'd54:begin
	fifo_WVALID_row[9][0]<=1'd0;
    fifo_WVALID_row[9][1]<=1'd0;
    fifo_WVALID_row[9][2]<=1'd0;
    fifo_WVALID_row[9][3]<=1'd0;	
	in_row[9][4]<=DO[7:0];
	in_row[9][5]<=DO[15:8];
	in_row[9][6]<=DO[23:16];
	in_row[9][7]<=DO[31:24];
	fifo_WVALID_row[9][4]<=1'd1;
    fifo_WVALID_row[9][5]<=1'd1;
    fifo_WVALID_row[9][6]<=1'd1;
    fifo_WVALID_row[9][7]<=1'd1;		
	end	
	7'd55:begin
	fifo_WVALID_row[9][4]<=1'd0;
    fifo_WVALID_row[9][5]<=1'd0;
    fifo_WVALID_row[9][6]<=1'd0;
    fifo_WVALID_row[9][7]<=1'd0;	
	in_row[10][0]<=DO[7:0];
	in_row[10][1]<=DO[15:8];
	in_row[10][2]<=DO[23:16];
	in_row[10][3]<=DO[31:24];
	fifo_WVALID_row[10][0]<=1'd1;
    fifo_WVALID_row[10][1]<=1'd1;
    fifo_WVALID_row[10][2]<=1'd1;
    fifo_WVALID_row[10][3]<=1'd1;		
	end	
	7'd56:begin
	fifo_WVALID_row[10][0]<=1'd0;
    fifo_WVALID_row[10][1]<=1'd0;
    fifo_WVALID_row[10][2]<=1'd0;
    fifo_WVALID_row[10][3]<=1'd0;	
	in_row[10][4]<=DO[7:0];
	in_row[10][5]<=DO[15:8];
	in_row[10][6]<=DO[23:16];
	in_row[10][7]<=DO[31:24];
	fifo_WVALID_row[10][4]<=1'd1;
    fifo_WVALID_row[10][5]<=1'd1;
    fifo_WVALID_row[10][6]<=1'd1;
    fifo_WVALID_row[10][7]<=1'd1;		
	end	
	7'd57:begin
	fifo_WVALID_row[10][4]<=1'd0;
    fifo_WVALID_row[10][5]<=1'd0;
    fifo_WVALID_row[10][6]<=1'd0;
    fifo_WVALID_row[10][7]<=1'd0;	
	in_row[11][0]<=DO[7:0];
	in_row[11][1]<=DO[15:8];
	in_row[11][2]<=DO[23:16];
	in_row[11][3]<=DO[31:24];	
	fifo_WVALID_row[11][0]<=1'd1;
    fifo_WVALID_row[11][1]<=1'd1;
    fifo_WVALID_row[11][2]<=1'd1;
    fifo_WVALID_row[11][3]<=1'd1;	
	end	
	7'd58:begin
	fifo_WVALID_row[11][0]<=1'd0;
    fifo_WVALID_row[11][1]<=1'd0;
    fifo_WVALID_row[11][2]<=1'd0;
    fifo_WVALID_row[11][3]<=1'd0;
	in_row[11][4]<=DO[7:0];
	in_row[11][5]<=DO[15:8];
	in_row[11][6]<=DO[23:16];
	in_row[11][7]<=DO[31:24];
	fifo_WVALID_row[11][4]<=1'd1;
    fifo_WVALID_row[11][5]<=1'd1;
    fifo_WVALID_row[11][6]<=1'd1;
    fifo_WVALID_row[11][7]<=1'd1;	
	end	
	7'd59:begin
	fifo_WVALID_row[11][4]<=1'd0;
    fifo_WVALID_row[11][5]<=1'd0;
    fifo_WVALID_row[11][6]<=1'd0;
    fifo_WVALID_row[11][7]<=1'd0;	
	in_row[12][0]<=DO[7:0];
	in_row[12][1]<=DO[15:8];
	in_row[12][2]<=DO[23:16];
	in_row[12][3]<=DO[31:24];
	fifo_WVALID_row[12][0]<=1'd1;
    fifo_WVALID_row[12][1]<=1'd1;
    fifo_WVALID_row[12][2]<=1'd1;
    fifo_WVALID_row[12][3]<=1'd1;		
	end	
	7'd60:begin
	fifo_WVALID_row[12][0]<=1'd0;
    fifo_WVALID_row[12][1]<=1'd0;
    fifo_WVALID_row[12][2]<=1'd0;
    fifo_WVALID_row[12][3]<=1'd0;	
	in_row[12][4]<=DO[7:0];
	in_row[12][5]<=DO[15:8];
	in_row[12][6]<=DO[23:16];
	in_row[12][7]<=DO[31:24];
	fifo_WVALID_row[12][4]<=1'd1;
    fifo_WVALID_row[12][5]<=1'd1;
    fifo_WVALID_row[12][6]<=1'd1;
    fifo_WVALID_row[12][7]<=1'd1;		
	end	
	7'd61:begin
	fifo_WVALID_row[12][4]<=1'd0;
    fifo_WVALID_row[12][5]<=1'd0;
    fifo_WVALID_row[12][6]<=1'd0;
    fifo_WVALID_row[12][7]<=1'd0;	
	in_row[13][0]<=DO[7:0];
	in_row[13][1]<=DO[15:8];
	in_row[13][2]<=DO[23:16];
	in_row[13][3]<=DO[31:24];	
	fifo_WVALID_row[13][0]<=1'd1;
    fifo_WVALID_row[13][1]<=1'd1;
    fifo_WVALID_row[13][2]<=1'd1;
    fifo_WVALID_row[13][3]<=1'd1;	
	end	
	7'd62:begin
	fifo_WVALID_row[13][0]<=1'd0;
    fifo_WVALID_row[13][1]<=1'd0;
    fifo_WVALID_row[13][2]<=1'd0;
    fifo_WVALID_row[13][3]<=1'd0;
	in_row[13][4]<=DO[7:0];
	in_row[13][5]<=DO[15:8];
	in_row[13][6]<=DO[23:16];
	in_row[13][7]<=DO[31:24];	
	fifo_WVALID_row[13][4]<=1'd1;
    fifo_WVALID_row[13][5]<=1'd1;
    fifo_WVALID_row[13][6]<=1'd1;
    fifo_WVALID_row[13][7]<=1'd1;
	end	
	7'd63:begin
	fifo_WVALID_row[13][4]<=1'd0;
    fifo_WVALID_row[13][5]<=1'd0;
    fifo_WVALID_row[13][6]<=1'd0;
    fifo_WVALID_row[13][7]<=1'd0;
	in_row[14][0]<=DO[7:0];
	in_row[14][1]<=DO[15:8];
	in_row[14][2]<=DO[23:16];
	in_row[14][3]<=DO[31:24];
	fifo_WVALID_row[14][0]<=1'd1;
    fifo_WVALID_row[14][1]<=1'd1;
    fifo_WVALID_row[14][2]<=1'd1;
    fifo_WVALID_row[14][3]<=1'd1;	
	end	
	7'd64:begin
	fifo_WVALID_row[14][0]<=1'd0;
    fifo_WVALID_row[14][1]<=1'd0;
    fifo_WVALID_row[14][2]<=1'd0;
    fifo_WVALID_row[14][3]<=1'd0;	
	in_row[14][4]<=DO[7:0];
	in_row[14][5]<=DO[15:8];
	in_row[14][6]<=DO[23:16];
	in_row[14][7]<=DO[31:24];
	fifo_WVALID_row[14][4]<=1'd1;
    fifo_WVALID_row[14][5]<=1'd1;
    fifo_WVALID_row[14][6]<=1'd1;
    fifo_WVALID_row[14][7]<=1'd1;		
	end		
	7'd65:begin
	fifo_WVALID_row[14][4]<=1'd0;
    fifo_WVALID_row[14][5]<=1'd0;
    fifo_WVALID_row[14][6]<=1'd0;
    fifo_WVALID_row[14][7]<=1'd0;	
	in_row[15][0]<=DO[7:0];
	in_row[15][1]<=DO[15:8];
	in_row[15][2]<=DO[23:16];
	in_row[15][3]<=DO[31:24];
	fifo_WVALID_row[15][0]<=1'd1;
    fifo_WVALID_row[15][1]<=1'd1;
    fifo_WVALID_row[15][2]<=1'd1;
    fifo_WVALID_row[15][3]<=1'd1;		
	end	
	7'd66:begin
	fifo_WVALID_row[15][0]<=1'd0;
    fifo_WVALID_row[15][1]<=1'd0;
    fifo_WVALID_row[15][2]<=1'd0;
    fifo_WVALID_row[15][3]<=1'd0;
	in_row[15][4]<=DO[7:0];
	in_row[15][5]<=DO[15:8];
	in_row[15][6]<=DO[23:16];
	in_row[15][7]<=DO[31:24];
	fifo_WVALID_row[15][4]<=1'd1;
    fifo_WVALID_row[15][5]<=1'd1;
    fifo_WVALID_row[15][6]<=1'd1;
    fifo_WVALID_row[15][7]<=1'd1;
	end
	7'd67:begin
	fifo_WVALID_row[15][4]<=1'd0;
    fifo_WVALID_row[15][5]<=1'd0;
    fifo_WVALID_row[15][6]<=1'd0;
    fifo_WVALID_row[15][7]<=1'd0;
	end
	//default:begin
	//in_row<=0;	
	//end
	endcase
//=============pointwise2============================================================		
end//always
















endmodule